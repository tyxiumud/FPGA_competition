module ds1302_module
(
    input CLK,
	 input RSTn,
	 
	 input [7:0]Start_Sig,
	 output Done_Sig,
	 
	 input [7:0]Time_Write_Data,
	 output [7:0]Time_Read_Data,
	 
	 output RST,
	 output SCLK,
	 inout SIO

);


	 
/***************************/
	 
wire [7:0]Words_Addr;
wire [7:0]Write_Data;
wire [1:0]Access_Start_Sig;
	 
wire [7:0]Read_Data;
wire Access_Done_Sig;
	 	 
cmd_control U1
(
	     .CLK( CLK ),
		  .RSTn( RSTn ),
		  .Start_Sig( Start_Sig ),               // �Ĵ�����д����/��ַ��input - from top
		  .Done_Sig( Done_Sig ),                 // �Ĵ�����д����źţ�output - to top
		  .Time_Write_Data( Time_Write_Data ),   // input - from top
		  .Time_Read_Data( Time_Read_Data ),     // output - to top
		  .Access_Done_Sig( Access_Done_Sig ),   // I2C��д����ź�: input - from U2
		  .Access_Start_Sig( Access_Start_Sig ), // ��д����: output - to U2
		  .Read_Data( Read_Data ),               // �����ļĴ�������: input - from U2         
		  .Words_Addr( Words_Addr ),             // �Ĵ����ĵ�ַ: output - to U2
		  .Write_Data( Write_Data )              // д��ļĴ���������: output - to U2
);
	 
	 /*****************************/
  
	 
i2c_com U2
(
	     .CLK( CLK ),
		  .RSTn( RSTn ),
		  .Start_Sig( Access_Start_Sig ),  // input - from  U1
		  .Words_Addr( Words_Addr ),       // input - from U1
		  .Write_Data( Write_Data ),       // input - from U1
		  .Read_Data( Read_Data ),         // output - to U1
		  .Done_Sig( Access_Done_Sig ),    // output - to U1
		  .RST( RST ),                     // DS1302��CE�źţ�output - to top
		  .SCLK( SCLK ),                   // DS1302��SCLK�źţ�output - to top
		  .SIO( SIO )                      // DS1302��SIO�źţ�output - to top
);
	 
	 /*****************************/
	 
endmodule
